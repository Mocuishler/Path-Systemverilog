module hello;
  initial 
    begin
      $display(signed'(1'h1-2'h2));;

    end
endmodule


